library verilog;
use verilog.vl_types.all;
entity division_vlg_vec_tst is
end division_vlg_vec_tst;
