library verilog;
use verilog.vl_types.all;
entity SignedVXL_vlg_sample_tst is
    port(
        A               : in     vl_logic_vector(31 downto 0);
        B               : in     vl_logic_vector(31 downto 0);
        CLK             : in     vl_logic;
        Start           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end SignedVXL_vlg_sample_tst;
