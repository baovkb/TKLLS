library verilog;
use verilog.vl_types.all;
entity SignedVXL_vlg_vec_tst is
end SignedVXL_vlg_vec_tst;
