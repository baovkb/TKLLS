library verilog;
use verilog.vl_types.all;
entity signedVXL_vlg_vec_tst is
end signedVXL_vlg_vec_tst;
